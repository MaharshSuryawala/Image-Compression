`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    22:11:16 11/01/2017 
// Design Name: 
// Module Name:    Multiplier_8x8 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Multiplier_8x8(
F00, F01, F02, F03, F04, F05, F06, F07,
F10, F11, F12, F13, F14, F15, F16, F17,
F20, F21, F22, F23, F24, F25, F26, F27,
F30, F31, F32, F33, F34, F35, F36, F37,
F40, F41, F42, F43, F44, F45, F46, F47,
F50, F51, F52, F53, F54, F55, F56, F57,
F60, F61, F62, F63, F64, F65, F66, F67,
F70, F71, F72, F73, F74, F75, F76, F77,

D00, D01, D02, D03, D04, D05, D06, D07,
D10, D11, D12, D13, D14, D15, D16, D17,
D20, D21, D22, D23, D24, D25, D26, D27,
D30, D31, D32, D33, D34, D35, D36, D37,
D40, D41, D42, D43, D44, D45, D46, D47,
D50, D51, D52, D53, D54, D55, D56, D57,
D60, D61, D62, D63, D64, D65, D66, D67,
D70, D71, D72, D73, D74, D75, D76, D77,

H00, H01, H02, H03, H04, H05, H06, H07,
H10, H11, H12, H13, H14, H15, H16, H17,
H20, H21, H22, H23, H24, H25, H26, H27,
H30, H31, H32, H33, H34, H35, H36, H37,
H40, H41, H42, H43, H44, H45, H46, H47,
H50, H51, H52, H53, H54, H55, H56, H57,
H60, H61, H62, H63, H64, H65, H66, H67,
H70, H71, H72, H73, H74, H75, H76, H77

);

/*input[15:0] H[7:0][7:0];
input[15:0] [7:0][7:0];
output[15:0] F[7:0][7:0];
*/

//D*H

output[15:0] F00, F01, F02, F03, F04, F05, F06, F07;
output[15:0] F10, F11, F12, F13, F14, F15, F16, F17;
output[15:0] F20, F21, F22, F23, F24, F25, F26, F27;
output[15:0] F30, F31, F32, F33, F34, F35, F36, F37;
output[15:0] F40, F41, F42, F43, F44, F45, F46, F47;
output[15:0] F50, F51, F52, F53, F54, F55, F56, F57;
output[15:0] F60, F61, F62, F63, F64, F65, F66, F67;
output[15:0] F70, F71, F72, F73, F74, F75, F76, F77;

wire[31:0] tF00, tF01, tF02, tF03, tF04, tF05, tF06, tF07;
wire[31:0] tF10, tF11, tF12, tF13, tF14, tF15, tF16, tF17;
wire[31:0] tF20, tF21, tF22, tF23, tF24, tF25, tF26, tF27;
wire[31:0] tF30, tF31, tF32, tF33, tF34, tF35, tF36, tF37;
wire[31:0] tF40, tF41, tF42, tF43, tF44, tF45, tF46, tF47;
wire[31:0] tF50, tF51, tF52, tF53, tF54, tF55, tF56, tF57;
wire[31:0] tF60, tF61, tF62, tF63, tF64, tF65, tF66, tF67;
wire[31:0] tF70, tF71, tF72, tF73, tF74, tF75, tF76, tF77;


input[15:0] D00, D01, D02, D03, D04, D05, D06, D07;
input[15:0] D10, D11, D12, D13, D14, D15, D16, D17;
input[15:0] D20, D21, D22, D23, D24, D25, D26, D27;
input[15:0] D30, D31, D32, D33, D34, D35, D36, D37;
input[15:0] D40, D41, D42, D43, D44, D45, D46, D47;
input[15:0] D50, D51, D52, D53, D54, D55, D56, D57;
input[15:0] D60, D61, D62, D63, D64, D65, D66, D67;
input[15:0] D70, D71, D72, D73, D74, D75, D76, D77;

input[15:0] H00, H01, H02, H03, H04, H05, H06, H07;
input[15:0] H10, H11, H12, H13, H14, H15, H16, H17;
input[15:0] H20, H21, H22, H23, H24, H25, H26, H27;
input[15:0] H30, H31, H32, H33, H34, H35, H36, H37;
input[15:0] H40, H41, H42, H43, H44, H45, H46, H47;
input[15:0] H50, H51, H52, H53, H54, H55, H56, H57;
input[15:0] H60, H61, H62, H63, H64, H65, H66, H67;
input[15:0] H70, H71, H72, H73, H74, H75, H76, H77;


assign tF00= D00*H00 + D01*H10 + D02*H20 + D03*H30 + D04*H40 + D05*H50 + D06*H60 + D07*H70; 
assign tF01= D00*H01 + D01*H11 + D02*H21 + D03*H31 + D04*H41 + D05*H51 + D06*H61 + D07*H71;
assign tF02= D00*H02 + D01*H12 + D02*H22 + D03*H32 + D04*H42 + D05*H52 + D06*H62 + D07*H72;
assign tF03= D00*H03 + D01*H13 + D02*H23 + D03*H33 + D04*H43 + D05*H53 + D06*H63 + D07*H73;
assign tF04= D00*H04 + D01*H14 + D02*H24 + D03*H34 + D04*H44 + D05*H54 + D06*H64 + D07*H74;
assign tF05= D00*H05 + D01*H15 + D02*H25 + D03*H35 + D04*H45 + D05*H55 + D06*H65 + D07*H75;
assign tF06= D00*H06 + D01*H16 + D02*H26 + D03*H36 + D04*H46 + D05*H56 + D06*H66 + D07*H76;
assign tF07= D00*H07 + D01*H17 + D02*H27 + D03*H37 + D04*H47 + D05*H57 + D06*H67 + D07*H77;

assign tF10= D10*H00 + D11*H10 + D12*H20 + D13*H30 + D14*H40 + D15*H50 + D16*H60 + D17*H70; 
assign tF11= D10*H01 + D11*H11 + D12*H21 + D13*H31 + D14*H41 + D15*H51 + D16*H61 + D17*H71;
assign tF12= D10*H02 + D11*H12 + D12*H22 + D13*H32 + D14*H42 + D15*H52 + D16*H62 + D17*H72;
assign tF13= D10*H03 + D11*H13 + D12*H23 + D13*H33 + D14*H43 + D15*H53 + D16*H63 + D17*H73;
assign tF14= D10*H04 + D11*H14 + D12*H24 + D13*H34 + D14*H44 + D15*H54 + D16*H64 + D17*H74;
assign tF15= D10*H05 + D11*H15 + D12*H25 + D13*H35 + D14*H45 + D15*H55 + D16*H65 + D17*H75;
assign tF16= D10*H06 + D11*H16 + D12*H26 + D13*H36 + D14*H46 + D15*H56 + D16*H66 + D17*H76;
assign tF17= D10*H07 + D11*H17 + D12*H27 + D13*H37 + D14*H47 + D15*H57 + D16*H67 + D17*H77;

assign tF20= D20*H00 + D21*H10 + D22*H20 + D23*H30 + D24*H40 + D25*H50 + D26*H60 + D27*H70; 
assign tF21= D20*H01 + D21*H11 + D22*H21 + D23*H31 + D24*H41 + D25*H51 + D26*H61 + D27*H71;
assign tF22= D20*H02 + D21*H12 + D22*H22 + D23*H32 + D24*H42 + D25*H52 + D26*H62 + D27*H72;
assign tF23= D20*H03 + D21*H13 + D22*H23 + D23*H33 + D24*H43 + D25*H53 + D26*H63 + D27*H73;
assign tF24= D20*H04 + D21*H14 + D22*H24 + D23*H34 + D24*H44 + D25*H54 + D26*H64 + D27*H74;
assign tF25= D20*H05 + D21*H15 + D22*H25 + D23*H35 + D24*H45 + D25*H55 + D26*H65 + D27*H75;
assign tF26= D20*H06 + D21*H16 + D22*H26 + D23*H36 + D24*H46 + D25*H56 + D26*H66 + D27*H76;
assign tF27= D20*H07 + D21*H17 + D22*H27 + D23*H37 + D24*H47 + D25*H57 + D26*H67 + D27*H77;

assign tF30= D30*H00 + D31*H10 + D32*H20 + D33*H30 + D34*H40 + D35*H50 + D36*H60 + D37*H70; 
assign tF31= D30*H01 + D31*H11 + D32*H21 + D33*H31 + D34*H41 + D35*H51 + D36*H61 + D37*H71;
assign tF32= D30*H02 + D31*H12 + D32*H22 + D33*H32 + D34*H42 + D35*H52 + D36*H62 + D37*H72;
assign tF33= D30*H03 + D31*H13 + D32*H23 + D33*H33 + D34*H43 + D35*H53 + D36*H63 + D37*H73;
assign tF34= D30*H04 + D31*H14 + D32*H24 + D33*H34 + D34*H44 + D35*H54 + D36*H64 + D37*H74;
assign tF35= D30*H05 + D31*H15 + D32*H25 + D33*H35 + D34*H45 + D35*H55 + D36*H65 + D37*H75;
assign tF36= D30*H06 + D31*H16 + D32*H26 + D33*H36 + D34*H46 + D35*H56 + D36*H66 + D37*H76;
assign tF37= D30*H07 + D31*H17 + D32*H27 + D33*H37 + D34*H47 + D35*H57 + D36*H67 + D37*H77;

assign tF40= D40*H00 + D41*H10 + D42*H20 + D43*H30 + D44*H40 + D45*H50 + D46*H60 + D47*H70; 
assign tF41= D40*H01 + D41*H11 + D42*H21 + D43*H31 + D44*H41 + D45*H51 + D46*H61 + D47*H71;
assign tF42= D40*H02 + D41*H12 + D42*H22 + D43*H32 + D44*H42 + D45*H52 + D46*H62 + D47*H72;
assign tF43= D40*H03 + D41*H13 + D42*H23 + D43*H33 + D44*H43 + D45*H53 + D46*H63 + D47*H73;
assign tF44= D40*H04 + D41*H14 + D42*H24 + D43*H34 + D44*H44 + D45*H54 + D46*H64 + D47*H74;
assign tF45= D40*H05 + D41*H15 + D42*H25 + D43*H35 + D44*H45 + D45*H55 + D46*H65 + D47*H75;
assign tF46= D40*H06 + D41*H16 + D42*H26 + D43*H36 + D44*H46 + D45*H56 + D46*H66 + D47*H76;
assign tF47= D40*H07 + D41*H17 + D42*H27 + D43*H37 + D44*H47 + D45*H57 + D46*H67 + D47*H77;

assign tF50= D50*H00 + D51*H10 + D52*H20 + D53*H30 + D54*H40 + D55*H50 + D56*H60 + D57*H70; 
assign tF51= D50*H01 + D51*H11 + D52*H21 + D53*H31 + D54*H41 + D55*H51 + D56*H61 + D57*H71;
assign tF52= D50*H02 + D51*H12 + D52*H22 + D53*H32 + D54*H42 + D55*H52 + D56*H62 + D57*H72;
assign tF53= D50*H03 + D51*H13 + D52*H23 + D53*H33 + D54*H43 + D55*H53 + D56*H63 + D57*H73;
assign tF54= D50*H04 + D51*H14 + D52*H24 + D53*H34 + D54*H44 + D55*H54 + D56*H64 + D57*H74;
assign tF55= D50*H05 + D51*H15 + D52*H25 + D53*H35 + D54*H45 + D55*H55 + D56*H65 + D57*H75;
assign tF56= D50*H06 + D51*H16 + D52*H26 + D53*H36 + D54*H46 + D55*H56 + D56*H66 + D57*H76;
assign tF57= D50*H07 + D51*H17 + D52*H27 + D53*H37 + D54*H47 + D55*H57 + D56*H67 + D57*H77;

assign tF60= D60*H00 + D61*H10 + D62*H20 + D63*H30 + D64*H40 + D65*H50 + D66*H60 + D67*H70; 
assign tF61= D60*H01 + D61*H11 + D62*H21 + D63*H31 + D64*H41 + D65*H51 + D66*H61 + D67*H71;
assign tF62= D60*H02 + D61*H12 + D62*H22 + D63*H32 + D64*H42 + D65*H52 + D66*H62 + D67*H72;
assign tF63= D60*H03 + D61*H13 + D62*H23 + D63*H33 + D64*H43 + D65*H53 + D66*H63 + D67*H73;
assign tF64= D60*H04 + D61*H14 + D62*H24 + D63*H34 + D64*H44 + D65*H54 + D66*H64 + D67*H74;
assign tF65= D60*H05 + D61*H15 + D62*H25 + D63*H35 + D64*H45 + D65*H55 + D66*H65 + D67*H75;
assign tF66= D60*H06 + D61*H16 + D62*H26 + D63*H36 + D64*H46 + D65*H56 + D66*H66 + D67*H76;
assign tF67= D60*H07 + D61*H17 + D62*H27 + D63*H37 + D64*H47 + D65*H57 + D66*H67 + D67*H77;

assign tF70= D70*H00 + D71*H10 + D72*H20 + D73*H30 + D74*H40 + D75*H50 + D76*H60 + D77*H70; 
assign tF71= D70*H01 + D71*H11 + D72*H21 + D73*H31 + D74*H41 + D75*H51 + D76*H61 + D77*H71;
assign tF72= D70*H02 + D71*H12 + D72*H22 + D73*H32 + D74*H42 + D75*H52 + D76*H62 + D77*H72;
assign tF73= D70*H03 + D71*H13 + D72*H23 + D73*H33 + D74*H43 + D75*H53 + D76*H63 + D77*H73;
assign tF74= D70*H04 + D71*H14 + D72*H24 + D73*H34 + D74*H44 + D75*H54 + D76*H64 + D77*H74;
assign tF75= D70*H05 + D71*H15 + D72*H25 + D73*H35 + D74*H45 + D75*H55 + D76*H65 + D77*H75;
assign tF76= D70*H06 + D71*H16 + D72*H26 + D73*H36 + D74*H46 + D75*H56 + D76*H66 + D77*H76;
assign tF77= D70*H07 + D71*H17 + D72*H27 + D73*H37 + D74*H47 + D75*H57 + D76*H67 + D77*H77;




assign F00= tF00[23:8];
assign F01= tF01[23:8];
assign F02= tF02[23:8];
assign F03= tF03[23:8];
assign F04= tF04[23:8];
assign F05= tF05[23:8];
assign F06= tF06[23:8];
assign F07= tF07[23:8];

assign F10= tF10[23:8];
assign F11= tF11[23:8];
assign F12= tF12[23:8];
assign F13= tF13[23:8];
assign F14= tF14[23:8];
assign F15= tF15[23:8];
assign F16= tF16[23:8];
assign F17= tF17[23:8];

assign F20= tF20[23:8];
assign F21= tF21[23:8];
assign F22= tF22[23:8];
assign F23= tF23[23:8];
assign F24= tF24[23:8];
assign F25= tF25[23:8];
assign F26= tF26[23:8];
assign F27= tF27[23:8];

assign F30= tF30[23:8];
assign F31= tF31[23:8];
assign F32= tF32[23:8];
assign F33= tF33[23:8];
assign F34= tF34[23:8];
assign F35= tF35[23:8];
assign F36= tF36[23:8];
assign F37= tF37[23:8];

assign F40= tF40[23:8];
assign F41= tF41[23:8];
assign F42= tF42[23:8];
assign F43= tF43[23:8];
assign F44= tF44[23:8];
assign F45= tF45[23:8];
assign F46= tF46[23:8];
assign F47= tF47[23:8];

assign F50= tF50[23:8];
assign F51= tF51[23:8];
assign F52= tF52[23:8];
assign F53= tF53[23:8];
assign F54= tF54[23:8];
assign F55= tF55[23:8];
assign F56= tF56[23:8];
assign F57= tF57[23:8];

assign F60= tF60[23:8];
assign F61= tF61[23:8];
assign F62= tF62[23:8];
assign F63= tF63[23:8];
assign F64= tF64[23:8];
assign F65= tF65[23:8];
assign F66= tF66[23:8];
assign F67= tF67[23:8];

assign F70= tF70[23:8];
assign F71= tF71[23:8];
assign F72= tF72[23:8];
assign F73= tF73[23:8];
assign F74= tF74[23:8];
assign F75= tF75[23:8];
assign F76= tF76[23:8];
assign F77= tF77[23:8];


/*assign F[1][0]= D[1][0]*H[0][0] + D[1][1]*H[1][0] + D[1][2]*H[2][0] + D[1][3]*H[3][0] + D[1][4]*H[4][0] + D[1][5]*H[5][0] + D[1][6]*H[6][0] + D[1][7]*H[7][0]; 
assign F[1][1]= D[1][0]*H[0][1] + D[1][1]*H[1][1] + D[1][2]*H[2][1] + D[1][3]*H[3][1] + D[1][4]*H[4][1] + D[1][5]*H[5][1] + D[1][6]*H[6][1] + D[1][7]*H[7][1];
assign F[1][2]= D[1][0]*H[0][2] + D[1][1]*H[1][2] + D[1][2]*H[2][2] + D[1][3]*H[3][2] + D[1][4]*H[4][2] + D[1][5]*H[5][2] + D[1][6]*H[6][2] + D[1][7]*H[7][2];
assign F[1][3]= D[1][0]*H[0][3] + D[1][1]*H[1][3] + D[1][2]*H[2][3] + D[1][3]*H[3][3] + D[1][4]*H[4][3] + D[1][5]*H[5][3] + D[1][6]*H[6][3] + D[1][7]*H[7][3];
assign F[1][4]= D[1][0]*H[0][4] + D[1][1]*H[1][4] + D[1][2]*H[2][4] + D[1][3]*H[3][4] + D[1][4]*H[4][4] + D[1][5]*H[5][4] + D[1][6]*H[6][4] + D[1][7]*H[7][4];
assign F[1][5]= D[1][0]*H[0][5] + D[1][1]*H[1][5] + D[1][2]*H[2][5] + D[1][3]*H[3][5] + D[1][4]*H[4][5] + D[1][5]*H[5][5] + D[1][6]*H[6][5] + D[1][7]*H[7][5];
assign F[1][6]= D[1][0]*H[0][6] + D[1][1]*H[1][6] + D[1][2]*H[2][6] + D[1][3]*H[3][6] + D[1][4]*H[4][6] + D[1][5]*H[5][6] + D[1][6]*H[6][6] + D[1][7]*H[7][6];
assign F[1][7]= D[1][0]*H[0][7] + D[1][1]*H[1][7] + D[1][2]*H[2][7] + D[1][3]*H[3][7] + D[1][4]*H[4][7] + D[1][5]*H[5][7] + D[1][6]*H[6][7] + D[1][7]*H[7][7];


assign F[2][0]= D[2][0]*H[0][0] + D[2][1]*H[1][0] + D[2][2]*H[2][0] + D[2][3]*H[3][0] + D[2][4]*H[4][0] + D[2][5]*H[5][0] + D[2][6]*H[6][0] + D[2][7]*H[7][0]; 
assign F[2][1]= D[2][0]*H[0][1] + D[2][1]*H[1][1] + D[2][2]*H[2][1] + D[2][3]*H[3][1] + D[2][4]*H[4][1] + D[2][5]*H[5][1] + D[2][6]*H[6][1] + D[2][7]*H[7][1];
assign F[2][2]= D[2][0]*H[0][2] + D[2][1]*H[1][2] + D[2][2]*H[2][2] + D[2][3]*H[3][2] + D[2][4]*H[4][2] + D[2][5]*H[5][2] + D[2][6]*H[6][2] + D[2][7]*H[7][2];
assign F[2][3]= D[2][0]*H[0][3] + D[2][1]*H[1][3] + D[2][2]*H[2][3] + D[2][3]*H[3][3] + D[2][4]*H[4][3] + D[2][5]*H[5][3] + D[2][6]*H[6][3] + D[2][7]*H[7][3];
assign F[2][4]= D[2][0]*H[0][4] + D[2][1]*H[1][4] + D[2][2]*H[2][4] + D[2][3]*H[3][4] + D[2][4]*H[4][4] + D[2][5]*H[5][4] + D[2][6]*H[6][4] + D[2][7]*H[7][4];
assign F[2][5]= D[2][0]*H[0][5] + D[2][1]*H[1][5] + D[2][2]*H[2][5] + D[2][3]*H[3][5] + D[2][4]*H[4][5] + D[2][5]*H[5][5] + D[2][6]*H[6][5] + D[2][7]*H[7][5];
assign F[2][6]= D[2][0]*H[0][6] + D[2][1]*H[1][6] + D[2][2]*H[2][6] + D[2][3]*H[3][6] + D[2][4]*H[4][6] + D[2][5]*H[5][6] + D[2][6]*H[6][6] + D[2][7]*H[7][6];
assign F[2][7]= D[2][0]*H[0][7] + D[2][1]*H[1][7] + D[2][2]*H[2][7] + D[2][3]*H[3][7] + D[2][4]*H[4][7] + D[2][5]*H[5][7] + D[2][6]*H[6][7] + D[2][7]*H[7][7];


assign F[3][0]= D[3][0]*H[0][0] + D[3][1]*H[1][0] + D[3][2]*H[2][0] + D[3][3]*H[3][0] + D[3][4]*H[4][0] + D[3][5]*H[5][0] + D[3][6]*H[6][0] + D[3][7]*H[7][0]; 
assign F[3][1]= D[3][0]*H[0][1] + D[3][1]*H[1][1] + D[3][2]*H[2][1] + D[3][3]*H[3][1] + D[3][4]*H[4][1] + D[3][5]*H[5][1] + D[3][6]*H[6][1] + D[3][7]*H[7][1];
assign F[3][2]= D[3][0]*H[0][2] + D[3][1]*H[1][2] + D[3][2]*H[2][2] + D[3][3]*H[3][2] + D[3][4]*H[4][2] + D[3][5]*H[5][2] + D[3][6]*H[6][2] + D[3][7]*H[7][2];
assign F[3][3]= D[3][0]*H[0][3] + D[3][1]*H[1][3] + D[3][2]*H[2][3] + D[3][3]*H[3][3] + D[3][4]*H[4][3] + D[3][5]*H[5][3] + D[3][6]*H[6][3] + D[3][7]*H[7][3];
assign F[3][4]= D[3][0]*H[0][4] + D[3][1]*H[1][4] + D[3][2]*H[2][4] + D[3][3]*H[3][4] + D[3][4]*H[4][4] + D[3][5]*H[5][4] + D[3][6]*H[6][4] + D[3][7]*H[7][4];
assign F[3][5]= D[3][0]*H[0][5] + D[3][1]*H[1][5] + D[3][2]*H[2][5] + D[3][3]*H[3][5] + D[3][4]*H[4][5] + D[3][5]*H[5][5] + D[3][6]*H[6][5] + D[3][7]*H[7][5];
assign F[3][6]= D[3][0]*H[0][6] + D[3][1]*H[1][6] + D[3][2]*H[2][6] + D[3][3]*H[3][6] + D[3][4]*H[4][6] + D[3][5]*H[5][6] + D[3][6]*H[6][6] + D[3][7]*H[7][6];
assign F[3][7]= D[3][0]*H[0][7] + D[3][1]*H[1][7] + D[3][2]*H[2][7] + D[3][3]*H[3][7] + D[3][4]*H[4][7] + D[3][5]*H[5][7] + D[3][6]*H[6][7] + D[3][7]*H[7][7];


assign F[4][0]= D[4][0]*H[0][0] + D[4][1]*H[1][0] + D[4][2]*H[2][0] + D[4][3]*H[3][0] + D[4][4]*H[4][0] + D[4][5]*H[5][0] + D[4][6]*H[6][0] + D[4][7]*H[7][0]; 
assign F[4][1]= D[4][0]*H[0][1] + D[4][1]*H[1][1] + D[4][2]*H[2][1] + D[4][3]*H[3][1] + D[4][4]*H[4][1] + D[4][5]*H[5][1] + D[4][6]*H[6][1] + D[4][7]*H[7][1];
assign F[4][2]= D[4][0]*H[0][2] + D[4][1]*H[1][2] + D[4][2]*H[2][2] + D[4][3]*H[3][2] + D[4][4]*H[4][2] + D[4][5]*H[5][2] + D[4][6]*H[6][2] + D[4][7]*H[7][2];
assign F[4][3]= D[4][0]*H[0][3] + D[4][1]*H[1][3] + D[4][2]*H[2][3] + D[4][3]*H[3][3] + D[4][4]*H[4][3] + D[4][5]*H[5][3] + D[4][6]*H[6][3] + D[4][7]*H[7][3];
assign F[4][4]= D[4][0]*H[0][4] + D[4][1]*H[1][4] + D[4][2]*H[2][4] + D[4][3]*H[3][4] + D[4][4]*H[4][4] + D[4][5]*H[5][4] + D[4][6]*H[6][4] + D[4][7]*H[7][4];
assign F[4][5]= D[4][0]*H[0][5] + D[4][1]*H[1][5] + D[4][2]*H[2][5] + D[4][3]*H[3][5] + D[4][4]*H[4][5] + D[4][5]*H[5][5] + D[4][6]*H[6][5] + D[4][7]*H[7][5];
assign F[4][6]= D[4][0]*H[0][6] + D[4][1]*H[1][6] + D[4][2]*H[2][6] + D[4][3]*H[3][6] + D[4][4]*H[4][6] + D[4][5]*H[5][6] + D[4][6]*H[6][6] + D[4][7]*H[7][6];
assign F[4][7]= D[4][0]*H[0][7] + D[4][1]*H[1][7] + D[4][2]*H[2][7] + D[4][3]*H[3][7] + D[4][4]*H[4][7] + D[4][5]*H[5][7] + D[4][6]*H[6][7] + D[4][7]*H[7][7];


assign F[5][0]= D[5][0]*H[0][0] + D[5][1]*H[1][0] + D[5][2]*H[2][0] + D[5][3]*H[3][0] + D[5][4]*H[4][0] + D[5][5]*H[5][0] + D[5][6]*H[6][0] + D[5][7]*H[7][0]; 
assign F[5][1]= D[5][0]*H[0][1] + D[5][1]*H[1][1] + D[5][2]*H[2][1] + D[5][3]*H[3][1] + D[5][4]*H[4][1] + D[5][5]*H[5][1] + D[5][6]*H[6][1] + D[5][7]*H[7][1];
assign F[5][2]= D[5][0]*H[0][2] + D[5][1]*H[1][2] + D[5][2]*H[2][2] + D[5][3]*H[3][2] + D[5][4]*H[4][2] + D[5][5]*H[5][2] + D[5][6]*H[6][2] + D[5][7]*H[7][2];
assign F[5][3]= D[5][0]*H[0][3] + D[5][1]*H[1][3] + D[5][2]*H[2][3] + D[5][3]*H[3][3] + D[5][4]*H[4][3] + D[5][5]*H[5][3] + D[5][6]*H[6][3] + D[5][7]*H[7][3];
assign F[5][4]= D[5][0]*H[0][4] + D[5][1]*H[1][4] + D[5][2]*H[2][4] + D[5][3]*H[3][4] + D[5][4]*H[4][4] + D[5][5]*H[5][4] + D[5][6]*H[6][4] + D[5][7]*H[7][4];
assign F[5][5]= D[5][0]*H[0][5] + D[5][1]*H[1][5] + D[5][2]*H[2][5] + D[5][3]*H[3][5] + D[5][4]*H[4][5] + D[5][5]*H[5][5] + D[5][6]*H[6][5] + D[5][7]*H[7][5];
assign F[5][6]= D[5][0]*H[0][6] + D[5][1]*H[1][6] + D[5][2]*H[2][6] + D[5][3]*H[3][6] + D[5][4]*H[4][6] + D[5][5]*H[5][6] + D[5][6]*H[6][6] + D[5][7]*H[7][6];
assign F[5][7]= D[5][0]*H[0][7] + D[5][1]*H[1][7] + D[5][2]*H[2][7] + D[5][3]*H[3][7] + D[5][4]*H[4][7] + D[5][5]*H[5][7] + D[5][6]*H[6][7] + D[5][7]*H[7][7];


assign F[6][0]= D[6][0]*H[0][0] + D[6][1]*H[1][0] + D[6][2]*H[2][0] + D[6][3]*H[3][0] + D[6][4]*H[4][0] + D[6][5]*H[5][0] + D[6][6]*H[6][0] + D[6][7]*H[7][0]; 
assign F[6][1]= D[6][0]*H[0][1] + D[6][1]*H[1][1] + D[6][2]*H[2][1] + D[6][3]*H[3][1] + D[6][4]*H[4][1] + D[6][5]*H[5][1] + D[6][6]*H[6][1] + D[6][7]*H[7][1];
assign F[6][2]= D[6][0]*H[0][2] + D[6][1]*H[1][2] + D[6][2]*H[2][2] + D[6][3]*H[3][2] + D[6][4]*H[4][2] + D[6][5]*H[5][2] + D[6][6]*H[6][2] + D[6][7]*H[7][2];
assign F[6][3]= D[6][0]*H[0][3] + D[6][1]*H[1][3] + D[6][2]*H[2][3] + D[6][3]*H[3][3] + D[6][4]*H[4][3] + D[6][5]*H[5][3] + D[6][6]*H[6][3] + D[6][7]*H[7][3];
assign F[6][4]= D[6][0]*H[0][4] + D[6][1]*H[1][4] + D[6][2]*H[2][4] + D[6][3]*H[3][4] + D[6][4]*H[4][4] + D[6][5]*H[5][4] + D[6][6]*H[6][4] + D[6][7]*H[7][4];
assign F[6][5]= D[6][0]*H[0][5] + D[6][1]*H[1][5] + D[6][2]*H[2][5] + D[6][3]*H[3][5] + D[6][4]*H[4][5] + D[6][5]*H[5][5] + D[6][6]*H[6][5] + D[6][7]*H[7][5];
assign F[6][6]= D[6][0]*H[0][6] + D[6][1]*H[1][6] + D[6][2]*H[2][6] + D[6][3]*H[3][6] + D[6][4]*H[4][6] + D[6][5]*H[5][6] + D[6][6]*H[6][6] + D[6][7]*H[7][6];
assign F[6][7]= D[6][0]*H[0][7] + D[6][1]*H[1][7] + D[6][2]*H[2][7] + D[6][3]*H[3][7] + D[6][4]*H[4][7] + D[6][5]*H[5][7] + D[6][6]*H[6][7] + D[6][7]*H[7][7];


assign F[7][0]= D[7][0]*H[0][0] + D[7][1]*H[1][0] + D[7][2]*H[2][0] + D[7][3]*H[3][0] + D[7][4]*H[4][0] + D[7][5]*H[5][0] + D[7][6]*H[6][0] + D[7][7]*H[7][0]; 
assign F[7][1]= D[7][0]*H[0][1] + D[7][1]*H[1][1] + D[7][2]*H[2][1] + D[7][3]*H[3][1] + D[7][4]*H[4][1] + D[7][5]*H[5][1] + D[7][6]*H[6][1] + D[7][7]*H[7][1];
assign F[7][2]= D[7][0]*H[0][2] + D[7][1]*H[1][2] + D[7][2]*H[2][2] + D[7][3]*H[3][2] + D[7][4]*H[4][2] + D[7][5]*H[5][2] + D[7][6]*H[6][2] + D[7][7]*H[7][2];
assign F[7][3]= D[7][0]*H[0][3] + D[7][1]*H[1][3] + D[7][2]*H[2][3] + D[7][3]*H[3][3] + D[7][4]*H[4][3] + D[7][5]*H[5][3] + D[7][6]*H[6][3] + D[7][7]*H[7][3];
assign F[7][4]= D[7][0]*H[0][4] + D[7][1]*H[1][4] + D[7][2]*H[2][4] + D[7][3]*H[3][4] + D[7][4]*H[4][4] + D[7][5]*H[5][4] + D[7][6]*H[6][4] + D[7][7]*H[7][4];
assign F[7][5]= D[7][0]*H[0][5] + D[7][1]*H[1][5] + D[7][2]*H[2][5] + D[7][3]*H[3][5] + D[7][4]*H[4][5] + D[7][5]*H[5][5] + D[7][6]*H[6][5] + D[7][7]*H[7][5];
assign F[7][6]= D[7][0]*H[0][6] + D[7][1]*H[1][6] + D[7][2]*H[2][6] + D[7][3]*H[3][6] + D[7][4]*H[4][6] + D[7][5]*H[5][6] + D[7][6]*H[6][6] + D[7][7]*H[7][6];
assign F[7][7]= D[7][0]*H[0][7] + D[7][1]*H[1][7] + D[7][2]*H[2][7] + D[7][3]*H[3][7] + D[7][4]*H[4][7] + D[7][5]*H[5][7] + D[7][6]*H[6][7] + D[7][7]*H[7][7];
*/

endmodule
